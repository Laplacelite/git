`timescale  1 ns / 1 ps
module ddr_master_top #(
    parameter ID_WIDTH                  = 4,
    parameter ADDR_WIDTH                = 32,
    parameter DATA_WIDTH                = 32,
    parameter AWUSER_WIDTH              = 1,
    parameter ARUSER_WIDTH              = 1, 
    parameter WUSER_WIDTH               = 1, 
    parameter RUSER_WIDTH               = 1,  
    parameter BUSER_WIDTH               = 1,
    parameter AW_LEN                    = 16,
    parameter AR_LEN                    = 16
)
(
        input   wire                                        m00_axi_init_axi_txn,
		output  wire                                        m00_axi_txn_done,
		output  wire                                        m00_axi_error,
		input   wire                                        m00_axi_aclk,
		input   wire                                        m00_axi_aresetn,
		output  wire        [C_M00_AXI_ID_WIDTH-1 : 0]      m00_axi_awid,
		output  wire        [C_M00_AXI_ADDR_WIDTH-1 : 0]    m00_axi_awaddr,
		output  wire        [7 : 0]                         m00_axi_awlen,
		output  wire        [2 : 0]                         m00_axi_awsize,
		output  wire        [1 : 0]                         m00_axi_awburst,
		output  wire                                        m00_axi_awlock,
		output  wire        [3 : 0]                         m00_axi_awcache,
		output  wire        [2 : 0]                         m00_axi_awprot,
		output  wire        [3 : 0]                         m00_axi_awqos,
		output  wire        [C_M00_AXI_AWUSER_WIDTH-1 : 0]  m00_axi_awuser,
		output  wire                                        m00_axi_awvalid,
		input   wire                                        m00_axi_awready,
		output  wire        [C_M00_AXI_DATA_WIDTH-1 : 0]    m00_axi_wdata,
		output  wire        [C_M00_AXI_DATA_WIDTH/8-1 : 0]  m00_axi_wstrb,
		output  wire                                        m00_axi_wlast,
		output  wire        [C_M00_AXI_WUSER_WIDTH-1 : 0]   m00_axi_wuser,
		output  wire                                        m00_axi_wvalid,
		input   wire                                        m00_axi_wready,
		input   wire        [C_M00_AXI_ID_WIDTH-1 : 0]      m00_axi_bid,
		input   wire        [1 : 0]                         m00_axi_bresp,
		input   wire        [C_M00_AXI_BUSER_WIDTH-1 : 0]   m00_axi_buser,
		input   wire                                        m00_axi_bvalid,
		output  wire                                        m00_axi_bready,
		output  wire        [C_M00_AXI_ID_WIDTH-1 : 0]      m00_axi_arid,
		output  wire        [C_M00_AXI_ADDR_WIDTH-1 : 0]    m00_axi_araddr,
		output  wire        [7 : 0]                         m00_axi_arlen,
		output  wire        [2 : 0]                         m00_axi_arsize,
		output  wire        [1 : 0]                         m00_axi_arburst,
		output  wire                                        m00_axi_arlock,
		output  wire        [3 : 0]                         m00_axi_arcache,
		output  wire        [2 : 0]                         m00_axi_arprot,
		output  wire        [3 : 0]                         m00_axi_arqos,
		output  wire        [C_M00_AXI_ARUSER_WIDTH-1 : 0]  m00_axi_aruser,
		output  wire                                        m00_axi_arvalid,
		input   wire                                        m00_axi_arready,
		input   wire        [C_M00_AXI_ID_WIDTH-1 : 0]      m00_axi_rid,
		input   wire        [C_M00_AXI_DATA_WIDTH-1 : 0]    m00_axi_rdata,
		input   wire        [1 : 0]                         m00_axi_rresp,
		input   wire                                        m00_axi_rlast,
		input   wire        [C_M00_AXI_RUSER_WIDTH-1 : 0]   m00_axi_ruser,
		input   wire                                        m00_axi_rvalid,
		output  wire                                        m00_axi_rready
	);

    ddr_master #(

    )
endmodule